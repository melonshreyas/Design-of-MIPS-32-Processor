module test_sub_adder();
sub_adder G1 (A,B,Diff);
reg [15:0] A,B;
wire [16:0] Sum;

initial
begin
$monitor ($time," Sum=%b, A=%b,B=%b", Sum, A,B);
end

initial
begin
#2  A=1174;B=40968;
#2  A=24105;B=18805;
#2  A=15294;B=42170;
#2  A=10660;B=62474;
#2  A=48898;B=60673;
#2  A=21376;B=17307;
#2  A=20382;B=6354;
#2  A=54944;B=56667;
#2  A=41745;B=52812;
#2  A=28900;B=44453;
#2  A=54507;B=33100;
#2  A=5989;B=12423;
#2  A=46515;B=45375;
#2  A=38493;B=40788;
#2  A=38237;B=15898;
#2  A=38254;B=48904;
#2  A=45643;B=44072;
#2  A=54047;B=44928;
#2  A=44079;B=21691;
#2  A=15312;B=27093;
#2  A=20616;B=31842;
#2  A=42183;B=29334;
#2  A=4135;B=55190;
#2  A=24750;B=40864;
#2  A=36559;B=63170;
end
