module alu_adder (A,B,Sum);
input [7:0] A,B;
output [8:0] Sum;
assign Sum=A+B;
endmodule
